`timescale 1ns / 1ps

module InstMem(Address, Instruction);
    input [31:0] Address;
    output reg [31:0] Instruction;

    always @(*)
        case (Address[9:2])
            8'd0: Instruction <= 32'h3c144000;
            8'd1: Instruction <= 32'h2294000c;
            8'd2: Instruction <= 32'h3c154000;
            8'd3: Instruction <= 32'h22b50010;
            8'd4: Instruction <= 32'h2010000f;
            8'd5: Instruction <= 32'h20110002;
            8'd6: Instruction <= 32'h20120200;
            8'd7: Instruction <= 32'h3c083332;
            8'd8: Instruction <= 32'h21083231;
            8'd9: Instruction <= 32'hae480000;
            8'd10: Instruction <= 32'h3c083136;
            8'd11: Instruction <= 32'h21083534;
            8'd12: Instruction <= 32'hae480004;
            8'd13: Instruction <= 32'h3c083231;
            8'd14: Instruction <= 32'h21083231;
            8'd15: Instruction <= 32'hae480008;
            8'd16: Instruction <= 32'h3c080036;
            8'd17: Instruction <= 32'h21083534;
            8'd18: Instruction <= 32'hae48000c;
            8'd19: Instruction <= 32'h20130400;
            8'd20: Instruction <= 32'h3c080000;
            8'd21: Instruction <= 32'h21083231;
            8'd22: Instruction <= 32'hae680000;
            8'd23: Instruction <= 32'h00102021;
            8'd24: Instruction <= 32'h00113021;
            8'd25: Instruction <= 32'h00122821;
            8'd26: Instruction <= 32'h00133821;
            8'd27: Instruction <= 32'h0c10006d;
            8'd28: Instruction <= 32'h20080000;
            8'd29: Instruction <= 32'h1048001e;
            8'd30: Instruction <= 32'h20080001;
            8'd31: Instruction <= 32'h1048001f;
            8'd32: Instruction <= 32'h20080002;
            8'd33: Instruction <= 32'h10480020;
            8'd34: Instruction <= 32'h20080003;
            8'd35: Instruction <= 32'h10480021;
            8'd36: Instruction <= 32'h20080004;
            8'd37: Instruction <= 32'h10480022;
            8'd38: Instruction <= 32'h20080005;
            8'd39: Instruction <= 32'h10480023;
            8'd40: Instruction <= 32'h20080006;
            8'd41: Instruction <= 32'h10480024;
            8'd42: Instruction <= 32'h20080007;
            8'd43: Instruction <= 32'h10480025;
            8'd44: Instruction <= 32'h20080008;
            8'd45: Instruction <= 32'h10480026;
            8'd46: Instruction <= 32'h20080009;
            8'd47: Instruction <= 32'h10480027;
            8'd48: Instruction <= 32'h2008000a;
            8'd49: Instruction <= 32'h10480028;
            8'd50: Instruction <= 32'h2008000b;
            8'd51: Instruction <= 32'h10480029;
            8'd52: Instruction <= 32'h2008000c;
            8'd53: Instruction <= 32'h1048002a;
            8'd54: Instruction <= 32'h2008000d;
            8'd55: Instruction <= 32'h1048002b;
            8'd56: Instruction <= 32'h2008000e;
            8'd57: Instruction <= 32'h1048002c;
            8'd58: Instruction <= 32'h2008000f;
            8'd59: Instruction <= 32'h1048002d;
            8'd60: Instruction <= 32'h2409013f;
            8'd61: Instruction <= 32'haea90000;
            8'd62: Instruction <= 32'h0810006c;
            8'd63: Instruction <= 32'h24090106;
            8'd64: Instruction <= 32'haea90000;
            8'd65: Instruction <= 32'h0810006c;
            8'd66: Instruction <= 32'h2409015b;
            8'd67: Instruction <= 32'haea90000;
            8'd68: Instruction <= 32'h0810006c;
            8'd69: Instruction <= 32'h2409014f;
            8'd70: Instruction <= 32'haea90000;
            8'd71: Instruction <= 32'h0810006c;
            8'd72: Instruction <= 32'h24090166;
            8'd73: Instruction <= 32'haea90000;
            8'd74: Instruction <= 32'h0810006c;
            8'd75: Instruction <= 32'h2409016d;
            8'd76: Instruction <= 32'haea90000;
            8'd77: Instruction <= 32'h0810006c;
            8'd78: Instruction <= 32'h2409017d;
            8'd79: Instruction <= 32'haea90000;
            8'd80: Instruction <= 32'h0810006c;
            8'd81: Instruction <= 32'h24090107;
            8'd82: Instruction <= 32'haea90000;
            8'd83: Instruction <= 32'h0810006c;
            8'd84: Instruction <= 32'h2409017f;
            8'd85: Instruction <= 32'haea90000;
            8'd86: Instruction <= 32'h0810006c;
            8'd87: Instruction <= 32'h2409016f;
            8'd88: Instruction <= 32'haea90000;
            8'd89: Instruction <= 32'h0810006c;
            8'd90: Instruction <= 32'h24090177;
            8'd91: Instruction <= 32'haea90000;
            8'd92: Instruction <= 32'h0810006c;
            8'd93: Instruction <= 32'h2409017c;
            8'd94: Instruction <= 32'haea90000;
            8'd95: Instruction <= 32'h0810006c;
            8'd96: Instruction <= 32'h24090139;
            8'd97: Instruction <= 32'haea90000;
            8'd98: Instruction <= 32'h0810006c;
            8'd99: Instruction <= 32'h2409015e;
            8'd100: Instruction <= 32'haea90000;
            8'd101: Instruction <= 32'h0810006c;
            8'd102: Instruction <= 32'h24090179;
            8'd103: Instruction <= 32'haea90000;
            8'd104: Instruction <= 32'h0810006c;
            8'd105: Instruction <= 32'h24090171;
            8'd106: Instruction <= 32'haea90000;
            8'd107: Instruction <= 32'h0810006c;
            8'd108: Instruction <= 32'h0810006c;
            8'd109: Instruction <= 32'h24020000;
            8'd110: Instruction <= 32'h00865022;
            8'd111: Instruction <= 32'h24080000;
            8'd112: Instruction <= 32'h0148082a;
            8'd113: Instruction <= 32'h1420000f;
            8'd114: Instruction <= 32'h24090000;
            8'd115: Instruction <= 32'h0126082a;
            8'd116: Instruction <= 32'h10200008;
            8'd117: Instruction <= 32'h01095820;
            8'd118: Instruction <= 32'h01655820;
            8'd119: Instruction <= 32'h816b0000;
            8'd120: Instruction <= 32'h01276020;
            8'd121: Instruction <= 32'h818c0000;
            8'd122: Instruction <= 32'h156c0002;
            8'd123: Instruction <= 32'h21290001;
            8'd124: Instruction <= 32'h08100073;
            8'd125: Instruction <= 32'h15260001;
            8'd126: Instruction <= 32'h20420001;
            8'd127: Instruction <= 32'h21080001;
            8'd128: Instruction <= 32'h08100070;
            8'd129: Instruction <= 32'h03e00008;
            default: Instruction <= 32'h00000000;
        endcase

endmodule